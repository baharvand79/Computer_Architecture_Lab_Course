module Adder(
	input [31:0] x0, x1,
	output [31:0] res
);
	assign res = x0 + x1;
endmodule 
module ARM();

endmodule
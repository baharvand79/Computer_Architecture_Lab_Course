module ID_Stage();
    input
endmodule